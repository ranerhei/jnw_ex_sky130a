magic
tech sky130A
magscale 1 2
timestamp 1737983866
<< locali >>
rect 585 3380 779 6437
rect 582 2754 779 3380
rect 585 2147 779 2754
rect 1734 5442 1926 7096
rect 1734 3826 1930 5442
rect 602 1998 702 2147
rect 1734 2096 1926 3826
rect 602 1908 976 1998
rect 1798 1998 1898 2096
rect 1156 1908 1898 1998
rect 602 1898 1898 1908
<< viali >>
rect 976 1908 1156 2088
<< metal1 >>
rect 1354 6912 1930 7104
rect 842 4876 906 6448
rect 970 6022 1162 6648
rect 1738 6050 1930 6912
rect 966 5706 1162 6022
rect 1354 5858 1930 6050
rect 966 5593 1158 5706
rect 836 4812 842 4876
rect 906 4812 912 4876
rect 842 2748 906 4812
rect 966 3653 1161 5593
rect 1428 4876 1492 4882
rect 1428 4806 1492 4812
rect 966 2444 1158 3653
rect 1738 3412 1930 5858
rect 1350 3220 1930 3412
rect 1738 3142 1930 3220
rect 1736 2914 1930 3142
rect 966 2232 1162 2444
rect 1736 2356 1928 2914
rect 970 2094 1162 2232
rect 1354 2164 1928 2356
rect 964 2088 1168 2094
rect 964 1908 976 2088
rect 1156 1908 1168 2088
rect 964 1902 1168 1908
<< via1 >>
rect 842 4812 906 4876
rect 1428 4812 1492 4876
<< metal2 >>
rect 842 4876 906 4882
rect 518 4812 842 4876
rect 906 4812 1428 4876
rect 1492 4812 1498 4876
rect 842 4806 906 4812
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 682 0 1 6344
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 682 0 1 2124
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 1 0 678 0 1 3180
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 682 0 1 4236
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1734044400
transform 1 0 682 0 1 5290
box -184 -128 1336 928
<< labels >>
flabel metal1 1504 3220 1696 3412 0 FreeSans 1600 0 0 0 IBNS_20U
port 0 nsew
flabel metal2 518 4812 582 4876 0 FreeSans 1600 0 0 0 IBPS_5U
port 2 nsew
flabel locali 1236 1898 1336 1998 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
<< end >>
